package gb_ppu_common_pkg;

// States for PPU Modes, Pixel FIFO, etc.

endpackage : gb_ppu_common_pkg

import gb_ppu_common_pkg::*;
/* Top Level Module for GameBoy PPU

Inputs:

Outputs:

*/
module gb_ppu();

endmodule : gb_ppu

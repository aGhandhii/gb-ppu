/* Top Level Testbench for PPU */
module gb_ppu_tb ();

endmodule : gb_ppu_tb
